module onewire_reset (
    input wire clk,
    input wire enable,
    output reg drive_low,
    output reg done
);
    // TODO
endmodule