module onewire_read (
    input wire clk,
    input wire enable,
    output reg drive_low,
    output reg [7:0] data_out,
    output reg done
);
    // TODO
endmodule